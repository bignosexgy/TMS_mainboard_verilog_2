//****************************************Copyright (c)***********************************//
//原子哥在线教学平台：www.yuanzige.com
//技术支持：www.openedv.com
//淘宝店铺：http://openedv.taobao.com 
//关注微信公众平台微信号："正点原子"，免费获取ZYNQ & FPGA & STM32 & LINUX资料。
//版权所有，盗版必究。
//Copyright(C) 正点原子 2018-2028
//All rights reserved	                               
//----------------------------------------------------------------------------------------
// File name:           uart_loop
// Last modified Date:  2019/10/8 17:25:36
// Last Version:        V1.1
// Descriptions:        串口数据环回模块
//----------------------------------------------------------------------------------------
// Created by:          正点原子
// Created date:        2019/10/8 17:25:36
// Version:             V1.0
// Descriptions:        The original version
//
//----------------------------------------------------------------------------------------
//****************************************************************************************//

module key_led_association(
    input	         	   sys_clk,                   //系统时钟
    input            	   sys_rst_n,                 //系统复位，低电平有效   
	
	input           [3:0]  key_push,
	output   reg    [3:0]  led_state 	
    );



//*****************************************************
//**                    main code
//*****************************************************


//reg define     
reg  [32:0] cnt_led;
reg  [1:0]  led_control;

//用于计数0.2s的计数器
always @ (posedge sys_clk or negedge sys_rst_n) begin
    if(!sys_rst_n)
        cnt_led<=24'd9_999_999;
    else if(cnt_led<24'd9_999_999)
        cnt_led<=cnt_led+1;
    else
        cnt_led<=0;
end 

//用于led灯状态的选择
always @(posedge sys_clk or negedge sys_rst_n) begin
    if (!sys_rst_n)
        led_control <= 2'b00;
    else if(cnt_led == 24'd9_999_999) 
        led_control <= led_control + 1'b1;
    else
        led_control <= led_control;
end

//识别按键，切换显示模式
always @(posedge sys_clk or negedge sys_rst_n) begin
    if(!sys_rst_n) begin
          led_state<=4'b 0000;
    end	
	else if(key_push[0]== 1)  //按键1按下时，从右向左的流水灯效果
        case (led_control)
            2'b00   : led_state<=4'b1000;
            2'b01   : led_state<=4'b0100;
            2'b10   : led_state<=4'b0010;
            2'b11   : led_state<=4'b0001;
            default  : led_state<=4'b0000;
        endcase
    else if (key_push[1]==1)  //按键2按下时，从左向右的流水灯效果
        case (led_control)
            2'b00   : led_state<=4'b0001;
            2'b01   : led_state<=4'b0010;
            2'b10   : led_state<=4'b0100;
            2'b11   : led_state<=4'b1000;
            default  : led_state<=4'b0000;
        endcase
    else if (key_push[2]==1)  //按键3按下时，LED闪烁
        case (led_control)
            2'b00   : led_state<=4'b1111;
            2'b01   : led_state<=4'b0000;
            2'b10   : led_state<=4'b1111;
            2'b11   : led_state<=4'b0000;
            default  : led_state<=4'b0000;
        endcase
    else if (key_push[3]==1)  //按键4按下时，LED全亮
        led_state=4'b1111;
    else
        led_state<=4'b0000;    //无按键按下时，LED熄灭  
	
end

endmodule 